// romtest.v

// Generated using ACDS version 13.0sp1 232 at 2016.11.22.07:06:40

`timescale 1 ps / 1 ps
module romtest (
		input  wire       clk_clk,              //      clk.clk
		input  wire       reset_reset_n,        //    reset.reset_n
		input  wire [7:0] rom_0_s1_address,     // rom_0_s1.address
		input  wire       rom_0_s1_debugaccess, //         .debugaccess
		input  wire       rom_0_s1_clken,       //         .clken
		input  wire       rom_0_s1_chipselect,  //         .chipselect
		input  wire       rom_0_s1_write,       //         .write
		output wire [7:0] rom_0_s1_readdata,    //         .readdata
		input  wire [7:0] rom_0_s1_writedata    //         .writedata
	);

	wire    rst_controller_reset_out_reset;     // rst_controller:reset_out -> rom_0:reset
	wire    rst_controller_reset_out_reset_req; // rst_controller:reset_req -> rom_0:reset_req

	romtest_rom_0 rom_0 (
		.clk         (clk_clk),                            //   clk1.clk
		.address     (rom_0_s1_address),                   //     s1.address
		.debugaccess (rom_0_s1_debugaccess),               //       .debugaccess
		.clken       (rom_0_s1_clken),                     //       .clken
		.chipselect  (rom_0_s1_chipselect),                //       .chipselect
		.write       (rom_0_s1_write),                     //       .write
		.readdata    (rom_0_s1_readdata),                  //       .readdata
		.writedata   (rom_0_s1_writedata),                 //       .writedata
		.reset       (rst_controller_reset_out_reset),     // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req)  //       .reset_req
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (1)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req  (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

endmodule
